//systemVerilog HDL for "ECE473", "sim_total_PDN_currentSinks_C4bumps_XL" "systemVerilog"


module sim_total_PDN_currentSinks_C4bumps_XL ( );

endmodule
