
--Create Entity:
--Library=ECE473,Cell=sim_total_PDN_currentSinks_C4bumps_XL,View=entity
--Time:Mon Jun 10 20:34:29 2024
--By:mlw375

LIBRARY ieee;
USE ieee.std_logic_1164.all;
ENTITY \sim_total_PDN_currentSinks_C4bumps_XL\ IS
END \sim_total_PDN_currentSinks_C4bumps_XL\;
